module moduleName (
  ports
  one 
  wo 
  thee
);
  
endmodule